grammar edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal Inst_t 'inst' lexer classes {Keyword, Reserved}, precedence=1;
