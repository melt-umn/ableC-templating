grammar edu:umn:cs:melt:exts:ableC:templating:concretesyntax;

--imports silver:langutil;

--imports edu:umn:cs:melt:ableC:concretesyntax;
--imports edu:umn:cs:melt:ableC:concretesyntax:lexerHack as lh;

imports edu:umn:cs:melt:ableC:abstractsyntax:host as ast;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction as ast;

exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateStructForwardDecl;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateStructDecl;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateFunctionDecl;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:usingDecl;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationTypeExpr;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationExpr;

exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateKeyword;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateParameters;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:templateStructKeyword;
exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:maybeAttributes;
