grammar edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instantiationExpr;

imports silver:langutil only ast;

imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:concretesyntax;

imports edu:umn:cs:melt:exts:ableC:templating:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:templating:concretesyntax:instKeyword;

marking terminal TemplateIdentifier_t /[A-Za-z_\$][A-Za-z_0-9\$]*/ lexer classes {Cidentifier};
terminal TemplateLParen_t '(';

disambiguate TemplateLParen_t, LParen_t {
  pluck TemplateLParen_t;
}

concrete productions top::PrimaryExpr_c
| id::TemplateIdentifier_t '<' params::TypeNames_c '>'
  { top.ast = templateDirectRefExpr(name(id.lexeme, location=id.location), params.ast, location=top.location); }
| id::TemplateIdentifier_t '<' params::TypeNames_c '>' '(' a::ArgumentExprList_c ')'
  { top.ast = templateDirectCallExpr(name(id.lexeme, location=id.location), params.ast, foldExpr(a.ast), location=top.location); }
| id::TemplateIdentifier_t '<' params::TypeNames_c '>' '(' ')'
  { top.ast = templateDirectCallExpr(name(id.lexeme, location=id.location), params.ast, nilExpr(), location=top.location); }
| id::TemplateIdentifier_t '(' a::ArgumentExprList_c ')'
  { top.ast = templateInferredDirectCallExpr(name(id.lexeme, location=id.location), foldExpr(a.ast), location=top.location); }
| id::TemplateIdentifier_t '(' ')'
  { top.ast = templateInferredDirectCallExpr(name(id.lexeme, location=id.location), nilExpr(), location=top.location); }
  -- For use in silver-ableC
| 'inst' id::Identifier_c '<' params::TypeNames_c '>'
  { top.ast = templateDirectRefExpr(id.ast, params.ast, location=top.location); }
| 'inst' id::Identifier_c '<' params::TypeNames_c '>' '(' a::ArgumentExprList_c ')'
  { top.ast = templateDirectCallExpr(id.ast, params.ast, foldExpr(a.ast), location=top.location); }
| 'inst' id::Identifier_c '<' params::TypeNames_c '>' '(' ')'
  { top.ast = templateDirectCallExpr(id.ast, params.ast, nilExpr(), location=top.location); }
